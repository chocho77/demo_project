module main

fn main() {
	println('Hello World!')
    println('Variables')
	name := 'Bob'
    age := 20
    large_number := i64(9999999999)
    println(name) 
    println(age)
    println(large_number)

}
